module ZiMoAmplify(
	input [ 255 : 0 ] ZiMo ,
	output [ 511 : 0 ] ZiMo_amp ) ;
	
	assign ZiMo_amp[ 1 : 0 ] = { 2{ZiMo[ 0 ]} } ;
	assign ZiMo_amp[ 3 : 2 ] = { 2{ZiMo[ 1 ]} } ;
	assign ZiMo_amp[ 5 : 4 ] = { 2{ZiMo[ 2 ]} } ;
	assign ZiMo_amp[ 7 : 6 ] = { 2{ZiMo[ 3 ]} } ;
	assign ZiMo_amp[ 9 : 8 ] = { 2{ZiMo[ 4 ]} } ;
	assign ZiMo_amp[ 11 : 10 ] = { 2{ZiMo[ 5 ]} } ;
	assign ZiMo_amp[ 13 : 12 ] = { 2{ZiMo[ 6 ]} } ;
	assign ZiMo_amp[ 15 : 14 ] = { 2{ZiMo[ 7 ]} } ;
	assign ZiMo_amp[ 17 : 16 ] = { 2{ZiMo[ 8 ]} } ;
	assign ZiMo_amp[ 19 : 18 ] = { 2{ZiMo[ 9 ]} } ;
	assign ZiMo_amp[ 21 : 20 ] = { 2{ZiMo[ 10 ]} } ;
	assign ZiMo_amp[ 23 : 22 ] = { 2{ZiMo[ 11 ]} } ;
	assign ZiMo_amp[ 25 : 24 ] = { 2{ZiMo[ 12 ]} } ;
	assign ZiMo_amp[ 27 : 26 ] = { 2{ZiMo[ 13 ]} } ;
	assign ZiMo_amp[ 29 : 28 ] = { 2{ZiMo[ 14 ]} } ;
	assign ZiMo_amp[ 31 : 30 ] = { 2{ZiMo[ 15 ]} } ;
	assign ZiMo_amp[ 33 : 32 ] = { 2{ZiMo[ 16 ]} } ;
	assign ZiMo_amp[ 35 : 34 ] = { 2{ZiMo[ 17 ]} } ;
	assign ZiMo_amp[ 37 : 36 ] = { 2{ZiMo[ 18 ]} } ;
	assign ZiMo_amp[ 39 : 38 ] = { 2{ZiMo[ 19 ]} } ;
	assign ZiMo_amp[ 41 : 40 ] = { 2{ZiMo[ 20 ]} } ;
	assign ZiMo_amp[ 43 : 42 ] = { 2{ZiMo[ 21 ]} } ;
	assign ZiMo_amp[ 45 : 44 ] = { 2{ZiMo[ 22 ]} } ;
	assign ZiMo_amp[ 47 : 46 ] = { 2{ZiMo[ 23 ]} } ;
	assign ZiMo_amp[ 49 : 48 ] = { 2{ZiMo[ 24 ]} } ;
	assign ZiMo_amp[ 51 : 50 ] = { 2{ZiMo[ 25 ]} } ;
	assign ZiMo_amp[ 53 : 52 ] = { 2{ZiMo[ 26 ]} } ;
	assign ZiMo_amp[ 55 : 54 ] = { 2{ZiMo[ 27 ]} } ;
	assign ZiMo_amp[ 57 : 56 ] = { 2{ZiMo[ 28 ]} } ;
	assign ZiMo_amp[ 59 : 58 ] = { 2{ZiMo[ 29 ]} } ;
	assign ZiMo_amp[ 61 : 60 ] = { 2{ZiMo[ 30 ]} } ;
	assign ZiMo_amp[ 63 : 62 ] = { 2{ZiMo[ 31 ]} } ;
	assign ZiMo_amp[ 65 : 64 ] = { 2{ZiMo[ 32 ]} } ;
	assign ZiMo_amp[ 67 : 66 ] = { 2{ZiMo[ 33 ]} } ;
	assign ZiMo_amp[ 69 : 68 ] = { 2{ZiMo[ 34 ]} } ;
	assign ZiMo_amp[ 71 : 70 ] = { 2{ZiMo[ 35 ]} } ;
	assign ZiMo_amp[ 73 : 72 ] = { 2{ZiMo[ 36 ]} } ;
	assign ZiMo_amp[ 75 : 74 ] = { 2{ZiMo[ 37 ]} } ;
	assign ZiMo_amp[ 77 : 76 ] = { 2{ZiMo[ 38 ]} } ;
	assign ZiMo_amp[ 79 : 78 ] = { 2{ZiMo[ 39 ]} } ;
	assign ZiMo_amp[ 81 : 80 ] = { 2{ZiMo[ 40 ]} } ;
	assign ZiMo_amp[ 83 : 82 ] = { 2{ZiMo[ 41 ]} } ;
	assign ZiMo_amp[ 85 : 84 ] = { 2{ZiMo[ 42 ]} } ;
	assign ZiMo_amp[ 87 : 86 ] = { 2{ZiMo[ 43 ]} } ;
	assign ZiMo_amp[ 89 : 88 ] = { 2{ZiMo[ 44 ]} } ;
	assign ZiMo_amp[ 91 : 90 ] = { 2{ZiMo[ 45 ]} } ;
	assign ZiMo_amp[ 93 : 92 ] = { 2{ZiMo[ 46 ]} } ;
	assign ZiMo_amp[ 95 : 94 ] = { 2{ZiMo[ 47 ]} } ;
	assign ZiMo_amp[ 97 : 96 ] = { 2{ZiMo[ 48 ]} } ;
	assign ZiMo_amp[ 99 : 98 ] = { 2{ZiMo[ 49 ]} } ;
	assign ZiMo_amp[ 101 : 100 ] = { 2{ZiMo[ 50 ]} } ;
	assign ZiMo_amp[ 103 : 102 ] = { 2{ZiMo[ 51 ]} } ;
	assign ZiMo_amp[ 105 : 104 ] = { 2{ZiMo[ 52 ]} } ;
	assign ZiMo_amp[ 107 : 106 ] = { 2{ZiMo[ 53 ]} } ;
	assign ZiMo_amp[ 109 : 108 ] = { 2{ZiMo[ 54 ]} } ;
	assign ZiMo_amp[ 111 : 110 ] = { 2{ZiMo[ 55 ]} } ;
	assign ZiMo_amp[ 113 : 112 ] = { 2{ZiMo[ 56 ]} } ;
	assign ZiMo_amp[ 115 : 114 ] = { 2{ZiMo[ 57 ]} } ;
	assign ZiMo_amp[ 117 : 116 ] = { 2{ZiMo[ 58 ]} } ;
	assign ZiMo_amp[ 119 : 118 ] = { 2{ZiMo[ 59 ]} } ;
	assign ZiMo_amp[ 121 : 120 ] = { 2{ZiMo[ 60 ]} } ;
	assign ZiMo_amp[ 123 : 122 ] = { 2{ZiMo[ 61 ]} } ;
	assign ZiMo_amp[ 125 : 124 ] = { 2{ZiMo[ 62 ]} } ;
	assign ZiMo_amp[ 127 : 126 ] = { 2{ZiMo[ 63 ]} } ;
	assign ZiMo_amp[ 129 : 128 ] = { 2{ZiMo[ 64 ]} } ;
	assign ZiMo_amp[ 131 : 130 ] = { 2{ZiMo[ 65 ]} } ;
	assign ZiMo_amp[ 133 : 132 ] = { 2{ZiMo[ 66 ]} } ;
	assign ZiMo_amp[ 135 : 134 ] = { 2{ZiMo[ 67 ]} } ;
	assign ZiMo_amp[ 137 : 136 ] = { 2{ZiMo[ 68 ]} } ;
	assign ZiMo_amp[ 139 : 138 ] = { 2{ZiMo[ 69 ]} } ;
	assign ZiMo_amp[ 141 : 140 ] = { 2{ZiMo[ 70 ]} } ;
	assign ZiMo_amp[ 143 : 142 ] = { 2{ZiMo[ 71 ]} } ;
	assign ZiMo_amp[ 145 : 144 ] = { 2{ZiMo[ 72 ]} } ;
	assign ZiMo_amp[ 147 : 146 ] = { 2{ZiMo[ 73 ]} } ;
	assign ZiMo_amp[ 149 : 148 ] = { 2{ZiMo[ 74 ]} } ;
	assign ZiMo_amp[ 151 : 150 ] = { 2{ZiMo[ 75 ]} } ;
	assign ZiMo_amp[ 153 : 152 ] = { 2{ZiMo[ 76 ]} } ;
	assign ZiMo_amp[ 155 : 154 ] = { 2{ZiMo[ 77 ]} } ;
	assign ZiMo_amp[ 157 : 156 ] = { 2{ZiMo[ 78 ]} } ;
	assign ZiMo_amp[ 159 : 158 ] = { 2{ZiMo[ 79 ]} } ;
	assign ZiMo_amp[ 161 : 160 ] = { 2{ZiMo[ 80 ]} } ;
	assign ZiMo_amp[ 163 : 162 ] = { 2{ZiMo[ 81 ]} } ;
	assign ZiMo_amp[ 165 : 164 ] = { 2{ZiMo[ 82 ]} } ;
	assign ZiMo_amp[ 167 : 166 ] = { 2{ZiMo[ 83 ]} } ;
	assign ZiMo_amp[ 169 : 168 ] = { 2{ZiMo[ 84 ]} } ;
	assign ZiMo_amp[ 171 : 170 ] = { 2{ZiMo[ 85 ]} } ;
	assign ZiMo_amp[ 173 : 172 ] = { 2{ZiMo[ 86 ]} } ;
	assign ZiMo_amp[ 175 : 174 ] = { 2{ZiMo[ 87 ]} } ;
	assign ZiMo_amp[ 177 : 176 ] = { 2{ZiMo[ 88 ]} } ;
	assign ZiMo_amp[ 179 : 178 ] = { 2{ZiMo[ 89 ]} } ;
	assign ZiMo_amp[ 181 : 180 ] = { 2{ZiMo[ 90 ]} } ;
	assign ZiMo_amp[ 183 : 182 ] = { 2{ZiMo[ 91 ]} } ;
	assign ZiMo_amp[ 185 : 184 ] = { 2{ZiMo[ 92 ]} } ;
	assign ZiMo_amp[ 187 : 186 ] = { 2{ZiMo[ 93 ]} } ;
	assign ZiMo_amp[ 189 : 188 ] = { 2{ZiMo[ 94 ]} } ;
	assign ZiMo_amp[ 191 : 190 ] = { 2{ZiMo[ 95 ]} } ;
	assign ZiMo_amp[ 193 : 192 ] = { 2{ZiMo[ 96 ]} } ;
	assign ZiMo_amp[ 195 : 194 ] = { 2{ZiMo[ 97 ]} } ;
	assign ZiMo_amp[ 197 : 196 ] = { 2{ZiMo[ 98 ]} } ;
	assign ZiMo_amp[ 199 : 198 ] = { 2{ZiMo[ 99 ]} } ;
	assign ZiMo_amp[ 201 : 200 ] = { 2{ZiMo[ 100 ]} } ;
	assign ZiMo_amp[ 203 : 202 ] = { 2{ZiMo[ 101 ]} } ;
	assign ZiMo_amp[ 205 : 204 ] = { 2{ZiMo[ 102 ]} } ;
	assign ZiMo_amp[ 207 : 206 ] = { 2{ZiMo[ 103 ]} } ;
	assign ZiMo_amp[ 209 : 208 ] = { 2{ZiMo[ 104 ]} } ;
	assign ZiMo_amp[ 211 : 210 ] = { 2{ZiMo[ 105 ]} } ;
	assign ZiMo_amp[ 213 : 212 ] = { 2{ZiMo[ 106 ]} } ;
	assign ZiMo_amp[ 215 : 214 ] = { 2{ZiMo[ 107 ]} } ;
	assign ZiMo_amp[ 217 : 216 ] = { 2{ZiMo[ 108 ]} } ;
	assign ZiMo_amp[ 219 : 218 ] = { 2{ZiMo[ 109 ]} } ;
	assign ZiMo_amp[ 221 : 220 ] = { 2{ZiMo[ 110 ]} } ;
	assign ZiMo_amp[ 223 : 222 ] = { 2{ZiMo[ 111 ]} } ;
	assign ZiMo_amp[ 225 : 224 ] = { 2{ZiMo[ 112 ]} } ;
	assign ZiMo_amp[ 227 : 226 ] = { 2{ZiMo[ 113 ]} } ;
	assign ZiMo_amp[ 229 : 228 ] = { 2{ZiMo[ 114 ]} } ;
	assign ZiMo_amp[ 231 : 230 ] = { 2{ZiMo[ 115 ]} } ;
	assign ZiMo_amp[ 233 : 232 ] = { 2{ZiMo[ 116 ]} } ;
	assign ZiMo_amp[ 235 : 234 ] = { 2{ZiMo[ 117 ]} } ;
	assign ZiMo_amp[ 237 : 236 ] = { 2{ZiMo[ 118 ]} } ;
	assign ZiMo_amp[ 239 : 238 ] = { 2{ZiMo[ 119 ]} } ;
	assign ZiMo_amp[ 241 : 240 ] = { 2{ZiMo[ 120 ]} } ;
	assign ZiMo_amp[ 243 : 242 ] = { 2{ZiMo[ 121 ]} } ;
	assign ZiMo_amp[ 245 : 244 ] = { 2{ZiMo[ 122 ]} } ;
	assign ZiMo_amp[ 247 : 246 ] = { 2{ZiMo[ 123 ]} } ;
	assign ZiMo_amp[ 249 : 248 ] = { 2{ZiMo[ 124 ]} } ;
	assign ZiMo_amp[ 251 : 250 ] = { 2{ZiMo[ 125 ]} } ;
	assign ZiMo_amp[ 253 : 252 ] = { 2{ZiMo[ 126 ]} } ;
	assign ZiMo_amp[ 255 : 254 ] = { 2{ZiMo[ 127 ]} } ;
	assign ZiMo_amp[ 257 : 256 ] = { 2{ZiMo[ 128 ]} } ;
	assign ZiMo_amp[ 259 : 258 ] = { 2{ZiMo[ 129 ]} } ;
	assign ZiMo_amp[ 261 : 260 ] = { 2{ZiMo[ 130 ]} } ;
	assign ZiMo_amp[ 263 : 262 ] = { 2{ZiMo[ 131 ]} } ;
	assign ZiMo_amp[ 265 : 264 ] = { 2{ZiMo[ 132 ]} } ;
	assign ZiMo_amp[ 267 : 266 ] = { 2{ZiMo[ 133 ]} } ;
	assign ZiMo_amp[ 269 : 268 ] = { 2{ZiMo[ 134 ]} } ;
	assign ZiMo_amp[ 271 : 270 ] = { 2{ZiMo[ 135 ]} } ;
	assign ZiMo_amp[ 273 : 272 ] = { 2{ZiMo[ 136 ]} } ;
	assign ZiMo_amp[ 275 : 274 ] = { 2{ZiMo[ 137 ]} } ;
	assign ZiMo_amp[ 277 : 276 ] = { 2{ZiMo[ 138 ]} } ;
	assign ZiMo_amp[ 279 : 278 ] = { 2{ZiMo[ 139 ]} } ;
	assign ZiMo_amp[ 281 : 280 ] = { 2{ZiMo[ 140 ]} } ;
	assign ZiMo_amp[ 283 : 282 ] = { 2{ZiMo[ 141 ]} } ;
	assign ZiMo_amp[ 285 : 284 ] = { 2{ZiMo[ 142 ]} } ;
	assign ZiMo_amp[ 287 : 286 ] = { 2{ZiMo[ 143 ]} } ;
	assign ZiMo_amp[ 289 : 288 ] = { 2{ZiMo[ 144 ]} } ;
	assign ZiMo_amp[ 291 : 290 ] = { 2{ZiMo[ 145 ]} } ;
	assign ZiMo_amp[ 293 : 292 ] = { 2{ZiMo[ 146 ]} } ;
	assign ZiMo_amp[ 295 : 294 ] = { 2{ZiMo[ 147 ]} } ;
	assign ZiMo_amp[ 297 : 296 ] = { 2{ZiMo[ 148 ]} } ;
	assign ZiMo_amp[ 299 : 298 ] = { 2{ZiMo[ 149 ]} } ;
	assign ZiMo_amp[ 301 : 300 ] = { 2{ZiMo[ 150 ]} } ;
	assign ZiMo_amp[ 303 : 302 ] = { 2{ZiMo[ 151 ]} } ;
	assign ZiMo_amp[ 305 : 304 ] = { 2{ZiMo[ 152 ]} } ;
	assign ZiMo_amp[ 307 : 306 ] = { 2{ZiMo[ 153 ]} } ;
	assign ZiMo_amp[ 309 : 308 ] = { 2{ZiMo[ 154 ]} } ;
	assign ZiMo_amp[ 311 : 310 ] = { 2{ZiMo[ 155 ]} } ;
	assign ZiMo_amp[ 313 : 312 ] = { 2{ZiMo[ 156 ]} } ;
	assign ZiMo_amp[ 315 : 314 ] = { 2{ZiMo[ 157 ]} } ;
	assign ZiMo_amp[ 317 : 316 ] = { 2{ZiMo[ 158 ]} } ;
	assign ZiMo_amp[ 319 : 318 ] = { 2{ZiMo[ 159 ]} } ;
	assign ZiMo_amp[ 321 : 320 ] = { 2{ZiMo[ 160 ]} } ;
	assign ZiMo_amp[ 323 : 322 ] = { 2{ZiMo[ 161 ]} } ;
	assign ZiMo_amp[ 325 : 324 ] = { 2{ZiMo[ 162 ]} } ;
	assign ZiMo_amp[ 327 : 326 ] = { 2{ZiMo[ 163 ]} } ;
	assign ZiMo_amp[ 329 : 328 ] = { 2{ZiMo[ 164 ]} } ;
	assign ZiMo_amp[ 331 : 330 ] = { 2{ZiMo[ 165 ]} } ;
	assign ZiMo_amp[ 333 : 332 ] = { 2{ZiMo[ 166 ]} } ;
	assign ZiMo_amp[ 335 : 334 ] = { 2{ZiMo[ 167 ]} } ;
	assign ZiMo_amp[ 337 : 336 ] = { 2{ZiMo[ 168 ]} } ;
	assign ZiMo_amp[ 339 : 338 ] = { 2{ZiMo[ 169 ]} } ;
	assign ZiMo_amp[ 341 : 340 ] = { 2{ZiMo[ 170 ]} } ;
	assign ZiMo_amp[ 343 : 342 ] = { 2{ZiMo[ 171 ]} } ;
	assign ZiMo_amp[ 345 : 344 ] = { 2{ZiMo[ 172 ]} } ;
	assign ZiMo_amp[ 347 : 346 ] = { 2{ZiMo[ 173 ]} } ;
	assign ZiMo_amp[ 349 : 348 ] = { 2{ZiMo[ 174 ]} } ;
	assign ZiMo_amp[ 351 : 350 ] = { 2{ZiMo[ 175 ]} } ;
	assign ZiMo_amp[ 353 : 352 ] = { 2{ZiMo[ 176 ]} } ;
	assign ZiMo_amp[ 355 : 354 ] = { 2{ZiMo[ 177 ]} } ;
	assign ZiMo_amp[ 357 : 356 ] = { 2{ZiMo[ 178 ]} } ;
	assign ZiMo_amp[ 359 : 358 ] = { 2{ZiMo[ 179 ]} } ;
	assign ZiMo_amp[ 361 : 360 ] = { 2{ZiMo[ 180 ]} } ;
	assign ZiMo_amp[ 363 : 362 ] = { 2{ZiMo[ 181 ]} } ;
	assign ZiMo_amp[ 365 : 364 ] = { 2{ZiMo[ 182 ]} } ;
	assign ZiMo_amp[ 367 : 366 ] = { 2{ZiMo[ 183 ]} } ;
	assign ZiMo_amp[ 369 : 368 ] = { 2{ZiMo[ 184 ]} } ;
	assign ZiMo_amp[ 371 : 370 ] = { 2{ZiMo[ 185 ]} } ;
	assign ZiMo_amp[ 373 : 372 ] = { 2{ZiMo[ 186 ]} } ;
	assign ZiMo_amp[ 375 : 374 ] = { 2{ZiMo[ 187 ]} } ;
	assign ZiMo_amp[ 377 : 376 ] = { 2{ZiMo[ 188 ]} } ;
	assign ZiMo_amp[ 379 : 378 ] = { 2{ZiMo[ 189 ]} } ;
	assign ZiMo_amp[ 381 : 380 ] = { 2{ZiMo[ 190 ]} } ;
	assign ZiMo_amp[ 383 : 382 ] = { 2{ZiMo[ 191 ]} } ;
	assign ZiMo_amp[ 385 : 384 ] = { 2{ZiMo[ 192 ]} } ;
	assign ZiMo_amp[ 387 : 386 ] = { 2{ZiMo[ 193 ]} } ;
	assign ZiMo_amp[ 389 : 388 ] = { 2{ZiMo[ 194 ]} } ;
	assign ZiMo_amp[ 391 : 390 ] = { 2{ZiMo[ 195 ]} } ;
	assign ZiMo_amp[ 393 : 392 ] = { 2{ZiMo[ 196 ]} } ;
	assign ZiMo_amp[ 395 : 394 ] = { 2{ZiMo[ 197 ]} } ;
	assign ZiMo_amp[ 397 : 396 ] = { 2{ZiMo[ 198 ]} } ;
	assign ZiMo_amp[ 399 : 398 ] = { 2{ZiMo[ 199 ]} } ;
	assign ZiMo_amp[ 401 : 400 ] = { 2{ZiMo[ 200 ]} } ;
	assign ZiMo_amp[ 403 : 402 ] = { 2{ZiMo[ 201 ]} } ;
	assign ZiMo_amp[ 405 : 404 ] = { 2{ZiMo[ 202 ]} } ;
	assign ZiMo_amp[ 407 : 406 ] = { 2{ZiMo[ 203 ]} } ;
	assign ZiMo_amp[ 409 : 408 ] = { 2{ZiMo[ 204 ]} } ;
	assign ZiMo_amp[ 411 : 410 ] = { 2{ZiMo[ 205 ]} } ;
	assign ZiMo_amp[ 413 : 412 ] = { 2{ZiMo[ 206 ]} } ;
	assign ZiMo_amp[ 415 : 414 ] = { 2{ZiMo[ 207 ]} } ;
	assign ZiMo_amp[ 417 : 416 ] = { 2{ZiMo[ 208 ]} } ;
	assign ZiMo_amp[ 419 : 418 ] = { 2{ZiMo[ 209 ]} } ;
	assign ZiMo_amp[ 421 : 420 ] = { 2{ZiMo[ 210 ]} } ;
	assign ZiMo_amp[ 423 : 422 ] = { 2{ZiMo[ 211 ]} } ;
	assign ZiMo_amp[ 425 : 424 ] = { 2{ZiMo[ 212 ]} } ;
	assign ZiMo_amp[ 427 : 426 ] = { 2{ZiMo[ 213 ]} } ;
	assign ZiMo_amp[ 429 : 428 ] = { 2{ZiMo[ 214 ]} } ;
	assign ZiMo_amp[ 431 : 430 ] = { 2{ZiMo[ 215 ]} } ;
	assign ZiMo_amp[ 433 : 432 ] = { 2{ZiMo[ 216 ]} } ;
	assign ZiMo_amp[ 435 : 434 ] = { 2{ZiMo[ 217 ]} } ;
	assign ZiMo_amp[ 437 : 436 ] = { 2{ZiMo[ 218 ]} } ;
	assign ZiMo_amp[ 439 : 438 ] = { 2{ZiMo[ 219 ]} } ;
	assign ZiMo_amp[ 441 : 440 ] = { 2{ZiMo[ 220 ]} } ;
	assign ZiMo_amp[ 443 : 442 ] = { 2{ZiMo[ 221 ]} } ;
	assign ZiMo_amp[ 445 : 444 ] = { 2{ZiMo[ 222 ]} } ;
	assign ZiMo_amp[ 447 : 446 ] = { 2{ZiMo[ 223 ]} } ;
	assign ZiMo_amp[ 449 : 448 ] = { 2{ZiMo[ 224 ]} } ;
	assign ZiMo_amp[ 451 : 450 ] = { 2{ZiMo[ 225 ]} } ;
	assign ZiMo_amp[ 453 : 452 ] = { 2{ZiMo[ 226 ]} } ;
	assign ZiMo_amp[ 455 : 454 ] = { 2{ZiMo[ 227 ]} } ;
	assign ZiMo_amp[ 457 : 456 ] = { 2{ZiMo[ 228 ]} } ;
	assign ZiMo_amp[ 459 : 458 ] = { 2{ZiMo[ 229 ]} } ;
	assign ZiMo_amp[ 461 : 460 ] = { 2{ZiMo[ 230 ]} } ;
	assign ZiMo_amp[ 463 : 462 ] = { 2{ZiMo[ 231 ]} } ;
	assign ZiMo_amp[ 465 : 464 ] = { 2{ZiMo[ 232 ]} } ;
	assign ZiMo_amp[ 467 : 466 ] = { 2{ZiMo[ 233 ]} } ;
	assign ZiMo_amp[ 469 : 468 ] = { 2{ZiMo[ 234 ]} } ;
	assign ZiMo_amp[ 471 : 470 ] = { 2{ZiMo[ 235 ]} } ;
	assign ZiMo_amp[ 473 : 472 ] = { 2{ZiMo[ 236 ]} } ;
	assign ZiMo_amp[ 475 : 474 ] = { 2{ZiMo[ 237 ]} } ;
	assign ZiMo_amp[ 477 : 476 ] = { 2{ZiMo[ 238 ]} } ;
	assign ZiMo_amp[ 479 : 478 ] = { 2{ZiMo[ 239 ]} } ;
	assign ZiMo_amp[ 481 : 480 ] = { 2{ZiMo[ 240 ]} } ;
	assign ZiMo_amp[ 483 : 482 ] = { 2{ZiMo[ 241 ]} } ;
	assign ZiMo_amp[ 485 : 484 ] = { 2{ZiMo[ 242 ]} } ;
	assign ZiMo_amp[ 487 : 486 ] = { 2{ZiMo[ 243 ]} } ;
	assign ZiMo_amp[ 489 : 488 ] = { 2{ZiMo[ 244 ]} } ;
	assign ZiMo_amp[ 491 : 490 ] = { 2{ZiMo[ 245 ]} } ;
	assign ZiMo_amp[ 493 : 492 ] = { 2{ZiMo[ 246 ]} } ;
	assign ZiMo_amp[ 495 : 494 ] = { 2{ZiMo[ 247 ]} } ;
	assign ZiMo_amp[ 497 : 496 ] = { 2{ZiMo[ 248 ]} } ;
	assign ZiMo_amp[ 499 : 498 ] = { 2{ZiMo[ 249 ]} } ;
	assign ZiMo_amp[ 501 : 500 ] = { 2{ZiMo[ 250 ]} } ;
	assign ZiMo_amp[ 503 : 502 ] = { 2{ZiMo[ 251 ]} } ;
	assign ZiMo_amp[ 505 : 504 ] = { 2{ZiMo[ 252 ]} } ;
	assign ZiMo_amp[ 507 : 506 ] = { 2{ZiMo[ 253 ]} } ;
	assign ZiMo_amp[ 509 : 508 ] = { 2{ZiMo[ 254 ]} } ;
	assign ZiMo_amp[ 511 : 510 ] = { 2{ZiMo[ 255 ]} } ;
	
endmodule